../wb_intercon/wb_intercon.vh